----------------------------------TILE 0 -----------------------------------------------  -- Y
("00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100", -- 1
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 1
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 2
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 2
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 3
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 3
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 4
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 4
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 5
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 5
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 6
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 6
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 7
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 7
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 8
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 8
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 9
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 9
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 10
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 10
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 11
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 11
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 12
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 12
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 13
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 13
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 14
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 14
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 15
"00011100","00011100","00011100","00011100","00011100","00011100","00011100","00011100",  -- 15
"11111100","11111100","11111100","11111100","11111100","11111100","11111100","11111100",  -- 16
"11111100","11111100","11111100","11111100","11111100","11111100","11111100","11111100",  -- 16
----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 16
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 16
----------------------------------TILE 2 -----------------------------------------------  -- Y
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 1
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 1
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 2
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 2
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 3
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 3
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 4
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 4
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 5
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 5
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 6
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 6
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 7
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 7
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 8
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 8
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 9
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 9
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 10
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 10
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 11
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 11
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 12
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 12
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 13
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 13
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 14
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 14
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 15
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 15
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 16
"11100000","11100000","11100000","11100000","11100000","11100000","11100000","11100000",  -- 16
----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 16
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111"); -- 16
