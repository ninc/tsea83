library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lab is
    	Port ( clk,rst : in  STD_LOGIC;
           	vgaRed, vgaGreen : out  STD_LOGIC_VECTOR (2 downto 0);
           	vgaBlue : out  STD_LOGIC_VECTOR (2 downto 1);
           	ca,cb,cc,cd,ce,cf,cg,dp, Hsync,Vsync : out  STD_LOGIC;
           	an : out  STD_LOGIC_VECTOR (3 downto 0));
end lab;

architecture Behavioral of lab is

component leddriver
    	Port ( clk,rst : in  STD_LOGIC;
           	ca,cb,cc,cd,ce,cf,cg,dp : out  STD_LOGIC;
           	an : out  STD_LOGIC_VECTOR (3 downto 0);
           	ledvalue : in  STD_LOGIC_VECTOR (15 downto 0));
end component;

  --Jacob
signal color : std_logic_vector(7 downto 0) := "00000000";
signal color_next : std_logic_vector(7 downto 0) := "00000000";
subtype color_t is std_logic_vector(7 downto 0);
type tile_array is array (integer range 0 to 65535) of color_t;
signal xctr,yctr : std_logic_vector(9 downto 0) := "0000000000";
alias y_tileminne : std_logic_vector(3 downto 0) is yctr(3 downto 0);
alias x_tileminne : std_logic_vector(3 downto 0) is xctr(3 downto 0);
alias x_grafikminne : std_logic_vector(6 downto 0) is xctr(9 downto 3);
alias y_grafikminne : std_logic_vector(5 downto 0) is yctr(9 downto 4);
signal pos_tileminne : integer range 0 to 65535 := 0;
signal aktuell_tile : std_logic_vector(7 downto 0) := "00000000";
signal tileminne : tile_array :=
----------------------------------TILE 0 -----------------------------------------------  -- Y
("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000", -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 0
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 0
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 1
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 1
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 2
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 2
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 3
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 3
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 4
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 4
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 5
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 5
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 6
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 6
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 7
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 7
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 8
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 8
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 9
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 9
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 10
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 10
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 11
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 11
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 12
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 12
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 13
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 13
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 14
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 14
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 15
"00011111","00011111","00011111","00011111","00011111","00011111","00011111","00011111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 0 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 1 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 2 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 3 -----------------------------------------------  -- Y
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 0
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 1
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 2
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 3
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 4
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 5
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 6
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 7
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 8
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 9
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 10
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 11
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 12
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 13
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 14
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15
"00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",  -- 15

----------------------------------TILE 4 -----------------------------------------------  -- Y
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 0
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 1
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 2
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 3
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 4
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 5
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 6
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 7
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 8
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 9
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15

----------------------------------TILE 5 -----------------------------------------------  -- Y
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 0
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 1
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 2
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 3
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 4
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 5
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 6
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 7
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 8
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 9
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 11
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 12
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 13
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 14
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 15

----------------------------------TILE 6 -----------------------------------------------  -- Y
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 0
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 1
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 2
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 3
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 4
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 5
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 6
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 7
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 8
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 9
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 10
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 11
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 12
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 13
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 14
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 15

----------------------------------TILE 7 -----------------------------------------------  -- Y
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 0
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 0
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 1
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 1
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 2
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 2
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 3
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 3
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 4
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 4
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 5
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 5
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 6
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 6
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 7
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 7
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 8
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 8
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 9
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 9
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 10
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 10
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 11
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 11
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 12
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 12
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 13
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 13
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 14
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 14
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000",  -- 15
"11111000","11111000","11111000","11111000","11111000","11111000","11111000","11111000"); -- 15


signal pos_grafikminne : integer range 0 to 1199 := 0;
subtype tile_t is std_logic_vector(7 downto 0);
type grafik_array is array(integer range 0 to 1199) of tile_t;
signal grafikminne : grafik_array :=
------------------------------------------- Grafikminne 1 ----------------------------------------------------  -- Y
("00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001", -- 00
"00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001",  -- 00
"00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001",  -- 00
"00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001",  -- 00
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 01
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 01
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 01
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 01
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 02
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 02
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 02
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 02
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 03
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 03
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 03
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 03
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 04
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 04
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 04
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 04
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 05
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 05
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 05
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 05
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 06
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 06
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 06
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 06
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 07
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 07
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 07
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 07
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 08
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 08
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 08
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 08
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 09
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 09
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 09
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 09
---------------------------------------------------------------------------------------------------------------------
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011","00000011",  -- 10
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 11
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 12
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 13
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 14
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 15
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 16
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 16
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 16
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 16
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 17
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 17
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 17
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 17
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 18
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 18
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 18
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 18
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 19
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 19
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 19
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 19
---------------------------------------------------------------------------------------------------------------------
"00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010",  -- 20
"00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010",  -- 20
"00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010",  -- 20
"00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010","00000010",  -- 20
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 21
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 21
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 21
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 21
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 22
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 22
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 22
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 22
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 23
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 23
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 23
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 23
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 24
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 24
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 24
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 24
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 25
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 25
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 25
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 25
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 26
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 26
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 26
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 26
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 27
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 27
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 27
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 27
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 28
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 28
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 28
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",  -- 28
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 29
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 29
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111",  -- 29
"11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111","11111111"); -- 29



--Given kod
--signal xctr,yctr : std_logic_vector(9 downto 0) := "0000000000";
alias rad : std_logic_vector(6 downto 0) is yctr(9 downto 3); -- i bildminnet
alias kol : std_logic_vector(6 downto 0) is xctr(9 downto 3);  -- i bildminnet
alias ypix : std_logic_vector(2 downto 0) is yctr(2 downto 0); -- i pixeln
alias xpix : std_logic_vector(2 downto 0) is xctr(2 downto 0);  -- i pixeln
signal pixel : std_logic_vector(1 downto 0) := "00";
signal a,b,c,d : std_logic_vector(0 to 79) := X"00000000000000000000";
signal a0,a1,a2,b0,b1,b2,c0,c1,c2 : std_logic := '0';
signal nr : std_logic_vector(3 downto 0) := "0000";
signal ctr : std_logic_vector(15 downto 0) := X"0000"; -- ?
signal hs : std_logic := '1';
signal vs : std_logic := '1';

begin 

--Pixel r�knare == 25MHz klocka till VGA
process(clk) begin
	if rising_edge(clk) then
		if rst='1' then
			pixel <= "00";
		else
			pixel <= pixel + 1;
       		end if;
     	end if;
end process;


-- Grafikminnet
process(clk) begin
	if rising_edge(clk) then
		if rst='1' then
			aktuell_tile <= "00000000";
		else		
			if y_grafikminne<30 and x_grafikminne<40 and pixel=0 then
				-- H�mta aktuell tile fr�n grafikminnet
				aktuell_tile <= grafikminne(pos_grafikminne);
			end if;
		end if;
	end if;
end process;

pos_grafikminne <= conv_integer(x_grafikminne) + 40*conv_integer(y_grafikminne);

--Tileminnet
process(clk) begin 
	if rising_edge(clk) then
		if y_grafikminne<30 and x_grafikminne<40 and pixel=1 then
			--L�gg in n�sta pixel fr�n aktuell rad
			color_next <= tileminne(pos_tileminne);
		end if;
	end if;
end process;

--R�kna ut n�sta position i tileminnet			
pos_tileminne <= 256*conv_integer(aktuell_tile) + 16*conv_integer(y_tileminne) + conv_integer(x_tileminne);
  
--Hsync
process(clk) begin
	if rising_edge(clk) then
      		if rst='1' then
         		xctr <= "0000000000";
      		elsif pixel=0 then
       			if xctr=799 then
         			xctr <= "0000000000";
       			else
         			xctr <= xctr + 1; -- Stega i X led			
       			end if;
      		end if;
      		-- 
      		if xctr=670 then
        		hs <= '0';
      		elsif xctr=766 then
        		hs <= '1';
      		end if;
    	end if;
end process;

-- Vsync
process(clk) begin
	if rising_edge(clk) then
      		if rst='1' then
        		yctr <= "0000000000";
      		elsif xctr=799 and pixel=0 then
       			if yctr=520 then
         			yctr <= "0000000000";
       			else
         			yctr <= yctr + 1; -- Stega i Y led
       			end if;
       			--
       			if yctr=490 then
         			vs <= '0';
       			elsif  yctr=491 then
         			vs <= '1';
       			end if;
      		end if;
    	end if;
end process;

-- S�tt Hsync, Vsync
Hsync <= hs;
Vsync <= vs;
  
-- VGA
process(clk) begin
    	if rising_edge(clk) then
      		if yctr<480 then
        		if xctr<640 then
          			if pixel=3 then
            				color <= color_next;
          			end if;
        		end if;
      		end if;
    	end if;
end process;

-- S�tt den nya f�rgen  
vgaRed(2 downto 0) <= color(7 downto 5);
vgaGreen(2 downto 0) <= color(4 downto 2);
vgaBlue(2 downto 1) <= color(1 downto 0);
  
  -- ************************************
  
process(clk) begin
     	if rising_edge(clk) then
       		if rst='1' then
         		ctr <= X"0000";
       		elsif yctr=0 and xctr=0 and pixel=0 then
         		ctr <= ctr+1;
       		end if;
     	end if;
end process;
       
  led: leddriver port map (clk,rst,ca,cb,cc,cd,ce,cf,cg,dp,an, ctr);
end Behavioral;

