library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lab is
    Port ( clk,rst : in  STD_LOGIC;
           vgaRed, vgaGreen : out  STD_LOGIC_VECTOR (2 downto 0);
           vgaBlue : out  STD_LOGIC_VECTOR (2 downto 1);
           ca,cb,cc,cd,ce,cf,cg,dp, Hsync,Vsync : out  STD_LOGIC;
           an : out  STD_LOGIC_VECTOR (3 downto 0));
end lab;

architecture Behavioral of lab is
  component leddriver
    Port ( clk,rst : in  STD_LOGIC;
           ca,cb,cc,cd,ce,cf,cg,dp : out  STD_LOGIC;
           an : out  STD_LOGIC_VECTOR (3 downto 0);
           ledvalue : in  STD_LOGIC_VECTOR (15 downto 0));
  end component;

  signal xctr,yctr : std_logic_vector(9 downto 0) := "0000000000";
  alias rad : std_logic_vector(6 downto 0) is yctr(9 downto 3); -- i bildminnet
  alias kol : std_logic_vector(6 downto 0) is xctr(9 downto 3);  -- i bildminnet
  alias ypix : std_logic_vector(2 downto 0) is yctr(2 downto 0); -- i pixeln
  alias xpix : std_logic_vector(2 downto 0) is xctr(2 downto 0);  -- i pixeln
  signal pixel : std_logic_vector(1 downto 0) := "00";
  signal a,b,c,d : std_logic_vector(0 to 79) := X"00000000000000000000";
  signal a0,a1,a2,b0,b1,b2,c0,c1,c2 : std_logic := '0';
  signal nr : std_logic_vector(3 downto 0) := "0000";
  signal ctr : std_logic_vector(15 downto 0) := X"0000";
  signal hs : std_logic := '1';
  signal vs : std_logic := '1';
  type ram_t is array (0 to 59) of std_logic_vector(0 to 79);

  constant glider : ram_t := ("00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000010000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000001010000000000000000000000000000000000000000000000000000",
                              "00000000000000011000000110000000000001100000000000000000000000000000000000000000",
                              "00000000000000100010000110000000000001100000000000000000000000000000000000000000",
                              "00011000000001000001000110000000000000000000000000000000000000000000000000000000",
                              "00011000000001000101100001010000000000000000000000000000000000000000000000000000",
                              "00000000000001000001000000010000000000000000000000000000000000000000000000000000",
                              "00000000000000100010000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000011000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000110000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000001000100000000000000000000000000000000000000000000000000000000",
                              "00000000000000000010000010000000100000000000000000000000000000000000000000000000",                     
                              "00000000110000000010001011000010100000000000000000000000000000000000000000000000",
                              "00000000110000000010000010001100000000000000000000000000000000000000000000000000",
                              "00000000000000000001000100001100000000000011000000000000000000000000000000000000",
                              "00000000000000000000110000001100000000000011000000000000000000000000000000000000",
                              "00000000000000000000000000000010100000000000000000000000000000000000000000000000",                     
                              "00000000000000000000000000000000100000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                              "00000000000000000000000000000000000000000000000000000000000000000000000000000000"
                              );
  signal bildminne : ram_t := glider;
  signal video : std_logic;
begin
  process(clk) begin
     if rising_edge(clk) then
       if rst='1' then
         pixel <= "00";
       else
         pixel <= pixel + 1;
       end if;
     end if;
  end process;


  process(clk) begin
    if rising_edge(clk) then
      if rst='1' then
         xctr <= "0000000000";
      elsif pixel=3 then
       if xctr=799 then
         xctr <= "0000000000";
       else
         xctr <= xctr + 1;
       end if;
      end if;
      -- 
      if xctr=670 then
        hs <= '0';
      elsif xctr=766 then
        hs <= '1';
      end if;
    end if;
  end process;

  process(clk) begin
    if rising_edge(clk) then
      if rst='1' then
        yctr <= "0000000000";
      elsif xctr=799 and pixel=0 then
       if yctr=520 then
         yctr <= "0000000000";
       else
         yctr <= yctr + 1;
       end if;
       --
       if yctr=490 then
         vs <= '0';
       elsif  yctr=491 then
         vs <= '1';
       end if;
      end if;
    end if;
  end process;
  Hsync <= hs;
  Vsync <= vs;

    -- bildminne
  process(clk) begin
    if rising_edge(clk) then
      if ypix=0 and xpix=0 and pixel=0 then
        if rad<60 then
          if kol=0 then
            a <= b;
            b <= c;
            if rad<59 then
              c <= bildminne(conv_integer(rad) + 1);     
            elsif rad=59 then
              c <= X"00000000000000000000";
            end if;
          elsif kol=80 then
            bildminne(conv_integer(rad)) <= d;     
          end if;     
        end if;
      end if;
    end if;
  end process;
  
  -- GoL
  process(clk) begin
    if rising_edge(clk) then
      if rad<60 and ypix=0 and xpix=0 then
        if pixel=1 then
          if kol < 79 then
            a2 <= a(conv_integer(kol+1));
            b2 <= b(conv_integer(kol+1));
            c2 <= c(conv_integer(kol+1));
          elsif kol=79 then
            a2 <= '0';
            b2 <= '0';
            c2 <= '0';
          end if;
          a0 <= a1; a1<=a2; 
          b0 <= b1; b1<=b2; 
          c0 <= c1; c1<=c2; 
        elsif pixel=2 then
          -- antal 1-or i omgivningen
          nr <= ("000" & a0) + ("000" & a1) + ("000" & a2) + ("000" & b0) + ("000" & b2) + ("000" & c0) + ("000" & c1) + ("000" & c2);
        elsif pixel=3 then
          if kol<80 then
            if nr=3 or (b1='1' and nr=2) then
              d(conv_integer(kol)) <= '1';
            else
              d(conv_integer(kol)) <= '0';
            end if;
          end if;
        end if;
      end if;
    end if;
  end process;

      
  -- video
  process(clk) begin
    if rising_edge(clk) then
      if yctr<480 then
        if xctr<640 then
          if pixel=3 then
            video <= b(conv_integer(kol));
          end if;
        end if;
      end if;
    end if;
  end process;
  
  vgaRed(2 downto 0) <= (video & video & video);
  vgaGreen(2 downto 0) <= (video & video & video);
  vgaBlue(2 downto 1) <= (video & video);
  
  -- ************************************
  
  process(clk) begin
     if rising_edge(clk) then
       if rst='1' then
         ctr <= X"0000";
       elsif yctr=0 and xctr=0 and pixel=0 then
         ctr <= ctr+1;
       end if;
     end if;
  end process;
       
  led: leddriver port map (clk,rst,ca,cb,cc,cd,ce,cf,cg,dp,an, ctr);
end Behavioral;

